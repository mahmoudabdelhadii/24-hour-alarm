module flashmemcont ()